<?xml version="1.0" encoding="UTF-8" standalone="yes"?>
<data>
    <accounts>
        <currency>
            <base>true</base>
            <code>RUB</code>
            <on>true</on>
            <rate>1.0</rate>
            <title>Ruble</title>
        </currency>
        <startAmount>5000.0</startAmount>
        <title>Wallet</title>
    </accounts>
    <accounts>
        <currency>
            <base>false</base>
            <code>USD</code>
            <on>true</on>
            <rate>1.5</rate>
            <title>Dollar</title>
        </currency>
        <startAmount>3500.0</startAmount>
        <title>Visa</title>
    </accounts>
    <accounts>
        <currency>
            <base>true</base>
            <code>RUB</code>
            <on>true</on>
            <rate>1.0</rate>
            <title>Ruble</title>
        </currency>
        <startAmount>1420.0</startAmount>
        <title>Deposit RUB</title>
    </accounts>
    <accounts>
        <currency>
            <base>false</base>
            <code>USD</code>
            <on>true</on>
            <rate>1.5</rate>
            <title>Dollar</title>
        </currency>
        <startAmount>2970.0</startAmount>
        <title>Deposit USD</title>
    </accounts>
    <articles>
        <title>Grocery</title>
    </articles>
    <articles>
        <title>Utilities</title>
    </articles>
    <articles>
        <title>Transport</title>
    </articles>
    <articles>
        <title>Interest rate</title>
    </articles>
    <currencies>
        <base>true</base>
        <code>RUB</code>
        <on>true</on>
        <rate>1.0</rate>
        <title>Ruble</title>
    </currencies>
    <currencies>
        <base>false</base>
        <code>USD</code>
        <on>true</on>
        <rate>1.5</rate>
        <title>Dollar</title>
    </currencies>
    <currencies>
        <base>false</base>
        <code>EUR</code>
        <on>true</on>
        <rate>2.4</rate>
        <title>Euro</title>
    </currencies>
    <currencies>
        <base>false</base>
        <code>UAH</code>
        <on>true</on>
        <rate>1.2</rate>
        <title>Hrivna</title>
    </currencies>
    <transactions>
        <account>
            <currency>
                <base>true</base>
                <code>RUB</code>
                <on>true</on>
                <rate>1.0</rate>
                <title>Ruble</title>
            </currency>
            <startAmount>1420.0</startAmount>
            <title>Deposit RUB</title>
        </account>
        <amount>-321.0</amount>
        <article>
            <title>Transport</title>
        </article>
        <date>2020-11-09T14:36:35.813Z</date>
        <notice>taxi</notice>
    </transactions>
    <transactions>
        <account>
            <currency>
                <base>false</base>
                <code>USD</code>
                <on>true</on>
                <rate>1.5</rate>
                <title>Dollar</title>
            </currency>
            <startAmount>3500.0</startAmount>
            <title>Visa</title>
        </account>
        <amount>-1000.0</amount>
        <article>
            <title>Utilities</title>
        </article>
        <date>2020-11-09T14:36:35.813Z</date>
        <notice>Second apt</notice>
    </transactions>
    <transactions>
        <account>
            <currency>
                <base>true</base>
                <code>RUB</code>
                <on>true</on>
                <rate>1.0</rate>
                <title>Ruble</title>
            </currency>
            <startAmount>5000.0</startAmount>
            <title>Wallet</title>
        </account>
        <amount>-812.0</amount>
        <article>
            <title>Grocery</title>
        </article>
        <date>2020-11-09T14:36:35.813Z</date>
        <notice>Eggs</notice>
    </transactions>
    <transactions>
        <account>
            <currency>
                <base>false</base>
                <code>USD</code>
                <on>true</on>
                <rate>1.5</rate>
                <title>Dollar</title>
            </currency>
            <startAmount>2970.0</startAmount>
            <title>Deposit USD</title>
        </account>
        <amount>136.0</amount>
        <article>
            <title>Interest rate</title>
        </article>
        <date>2020-01-14T14:36:35.813Z</date>
        <notice></notice>
    </transactions>
    <transfers>
        <date>2020-11-09T14:36:35.813Z</date>
        <fromAccount>
            <currency>
                <base>false</base>
                <code>USD</code>
                <on>true</on>
                <rate>1.5</rate>
                <title>Dollar</title>
            </currency>
            <startAmount>3500.0</startAmount>
            <title>Visa</title>
        </fromAccount>
        <fromAmount>250.0</fromAmount>
        <notice></notice>
        <toAccount>
            <currency>
                <base>true</base>
                <code>RUB</code>
                <on>true</on>
                <rate>1.0</rate>
                <title>Ruble</title>
            </currency>
            <startAmount>5000.0</startAmount>
            <title>Wallet</title>
        </toAccount>
        <toAmount>250.0</toAmount>
    </transfers>
    <transfers>
        <date>2020-11-09T14:36:35.813Z</date>
        <fromAccount>
            <currency>
                <base>false</base>
                <code>USD</code>
                <on>true</on>
                <rate>1.5</rate>
                <title>Dollar</title>
            </currency>
            <startAmount>2970.0</startAmount>
            <title>Deposit USD</title>
        </fromAccount>
        <fromAmount>192.0</fromAmount>
        <notice></notice>
        <toAccount>
            <currency>
                <base>true</base>
                <code>RUB</code>
                <on>true</on>
                <rate>1.0</rate>
                <title>Ruble</title>
            </currency>
            <startAmount>1420.0</startAmount>
            <title>Deposit RUB</title>
        </toAccount>
        <toAmount>192.0</toAmount>
    </transfers>
    <transfers>
        <date>2020-11-09T14:36:35.813Z</date>
        <fromAccount>
            <currency>
                <base>true</base>
                <code>RUB</code>
                <on>true</on>
                <rate>1.0</rate>
                <title>Ruble</title>
            </currency>
            <startAmount>5000.0</startAmount>
            <title>Wallet</title>
        </fromAccount>
        <fromAmount>576.0</fromAmount>
        <notice></notice>
        <toAccount>
            <currency>
                <base>false</base>
                <code>USD</code>
                <on>true</on>
                <rate>1.5</rate>
                <title>Dollar</title>
            </currency>
            <startAmount>2970.0</startAmount>
            <title>Deposit USD</title>
        </toAccount>
        <toAmount>557.0</toAmount>
    </transfers>
</data>
